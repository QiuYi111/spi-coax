`timescale 1ns / 1ps

`include "tb_common.vh"

module tb_cdr;

    // ========================================================================
    // Test Control
    // ========================================================================
    reg test_failed;
    integer check_count, pass_count, fail_count;
    string section_name;

    // ========================================================================
    // DUT Signals
    // ========================================================================
    reg clk_link;
    reg rst_n;
    reg manch_in;
    wire bit_out;
    wire bit_valid;
    wire locked;

    // ========================================================================
    // Clock Generation (200MHz)
    // ========================================================================
    parameter real CLK_PERIOD = 5.0;  // 200MHz
    
    initial begin
        clk_link = 0;
        forever #(CLK_PERIOD/2) clk_link = ~clk_link;
    end

    // ========================================================================
    // DUT Instantiation
    // ========================================================================
    cdr_4x_oversampling u_dut (
        .clk_link(clk_link),
        .rst_n(rst_n),
        .manch_in(manch_in),
        .bit_out(bit_out),
        .bit_valid(bit_valid),
        .locked(locked)
    );

    // ========================================================================
    // Manchester Stream Generator
    // ========================================================================
    
    // Generate Manchester bit (0 -> 01, 1 -> 10) at 50 Mbps
    task send_manchester_bit;
        input bit_val;
        input real jitter_percent;  // Optional jitter
        real half_bit_time;
        real actual_time;
        begin
            // 50 Mbps = 20ns bit period, 10ns per half-bit
            half_bit_time = 10.0;
            
            if (bit_val == 0) begin
                // Encode 0 as 01
                actual_time = add_jitter(half_bit_time, jitter_percent);
                manch_in = 0;
                #actual_time;
                actual_time = add_jitter(half_bit_time, jitter_percent);
                manch_in = 1;
                #actual_time;
            end else begin
                // Encode 1 as 10
                actual_time = add_jitter(half_bit_time, jitter_percent);
                manch_in = 1;
                #actual_time;
                actual_time = add_jitter(half_bit_time, jitter_percent);
                manch_in = 0;
                #actual_time;
            end
        end
    endtask
    
    // Send training sequence (alternating pattern for lock)
    task send_training_sequence;
        input integer num_bits;
        integer i;
        begin
            for (i = 0; i < num_bits; i = i + 1) begin
                send_manchester_bit(i % 2, 0.0);
            end
        end
    endtask
    
    // Send data pattern
    task send_data_pattern;
        input [31:0] data;
        input integer num_bits;
        integer i;
        begin
            for (i = num_bits-1; i >= 0; i = i - 1) begin
                send_manchester_bit(data[i], 0.0);
            end
        end
    endtask
    
    // Send with bit errors
    task send_with_errors;
        input bit_val;
        input integer error_rate_ppm;
        reg actual_bit;
        begin
            actual_bit = inject_bit_error(bit_val, error_rate_ppm);
            send_manchester_bit(actual_bit, 0.0);
        end
    endtask

    // ========================================================================
    // Monitoring and Verification
    // ========================================================================
    
    integer lock_time;
    integer bits_received;
    integer bits_expected;
    integer bit_errors;
    integer lock_count;
    integer unlock_count;
    
    // Monitor lock acquisition
    always @(posedge locked) begin
        lock_time = $time;
        lock_count = lock_count + 1;
        $display("[CDR LOCK] Acquired at time %0t (%.2f us)", lock_time, lock_time / 1000.0);
    end
    
    always @(negedge locked) begin
        unlock_count = unlock_count + 1;
        $display("[CDR UNLOCK] Lost lock at time %0t", $time);
    end
    
    // Count received bits
    always @(posedge clk_link) begin
        if (bit_valid) begin
            bits_received = bits_received + 1;
        end
    end
    
    // Verify received bits
    task verify_received_bits;
        input [31:0] expected_data;
        input integer num_bits;
        reg [31:0] received_data;
        integer i;
        integer timeout;
        begin
            received_data = 0;
            timeout = 0;
            
            for (i = num_bits-1; i >= 0; i = i - 1) begin
                // Wait for bit_valid
                timeout = 0;
                while (!bit_valid && timeout < 1000) begin
                    @(posedge clk_link);
                    timeout = timeout + 1;
                end
                
                if (timeout >= 1000) begin
                    $error("[VERIFY] Timeout waiting for bit %0d", i);
                    bit_errors = bit_errors + 1;
                end else begin
                    received_data[i] = bit_out;
                    @(posedge clk_link);
                end
            end
            
            // Check match
            if (received_data === expected_data) begin
                $display("[VERIFY] PASS: Received %h matches expected %h", received_data, expected_data);
            end else begin
                $error("[VERIFY] FAIL: Received %h, expected %h", received_data, expected_data);
                bit_errors = bit_errors + 1;
            end
        end
    endtask

    // ========================================================================
    // Test Scenarios
    // ========================================================================
    
    task reset_test;
        begin
            `TEST_SECTION("Reset and Initialization")
            
            rst_n = 0;
            manch_in = 0;
            
            #200;
            rst_n = 1;
            #100;
            
            `ASSERT(locked === 1'b0, "CDR should not be locked after reset")
            `ASSERT(bit_valid === 1'b0, "No valid bits should be output after reset")
            
            $display("Reset test completed");
        end
    endtask
    
    task lock_acquisition_test;
        integer start_time;
        integer lock_duration;
        begin
            `TEST_SECTION("Lock Acquisition")
            
            start_time = $time;
            
            // Send training sequence
            send_training_sequence(100);
            
            // Wait for lock
            wait(locked);
            
            lock_duration = $time - start_time;
            
            $display("[LOCK ACQUISITION] Time to lock: %0d ns (%.2f us)", 
                     lock_duration, lock_duration / 1000.0);
            
            // Should lock within reasonable time (typically < 1ms)
            `CHECK_RANGE(lock_duration, 0, 1000000, "Lock Acquisition Time (ns)")
            
            $display("Lock acquisition test completed");
        end
    endtask
    
    task data_recovery_test;
        reg [31:0] test_data;
        begin
            `TEST_SECTION("Data Recovery - Simple Pattern")
            
            // Ensure locked
            if (!locked) begin
                send_training_sequence(100);
                wait(locked);
            end
            
            // Send known data pattern
            test_data = 32'hA5A5A5A5;
            bits_expected = 32;
            
            $display("Sending data pattern: %h", test_data);
            send_data_pattern(test_data, 32);
            
            // Verify (note: need to collect bits separately in real implementation)
            // For now, just check we got valid bits
            `ASSERT(bits_received > 0, "Should have received some bits")
            
            $display("Data recovery test completed");
        end
    endtask
    
    task alternating_pattern_test;
        integer i;
        begin
            `TEST_SECTION("Alternating Bit Pattern")
            
            // Ensure locked
            if (!locked) begin
                send_training_sequence(50);
                wait(locked);
            end
            
            // Send alternating pattern
            for (i = 0; i < 32; i = i send_manchester_bit(i % 2, 0.0);
            end
            
            $display("Alternating pattern test completed");
        end
    endtask
    
    task all_zeros_test;
        integer i;
        begin
            `TEST_SECTION("All Zeros Pattern")
            
            if (!locked) begin
                send_training_sequence(50);
                wait(locked);
            end
            
            for (i = 0; i < 16; i = i + 1) begin
                send_manchester_bit(1'b0, 0.0);
            end
            
            $display("All zeros test completed");
        end
    endtask
    
    task all_ones_test;
        integer i;
        begin
            `TEST_SECTION("All Ones Pattern")
            
            if (!locked) begin
                send_training_sequence(50);
                wait(locked);
            end
            
            for (i = 0; i < 16; i = i + 1) begin
                send_manchester_bit(1'b1, 0.0);
            end
            
            $display("All ones test completed");
        end
    endtask
    
    task jitter_tolerance_test;
        integer i;
        real jitter_levels [0:3];
        integer j;
        begin
            `TEST_SECTION("Jitter Tolerance")
            
            // Test different jitter levels
            jitter_levels[0] = 0.0;   // No jitter
            jitter_levels[1] = 5.0;   // 5% jitter
            jitter_levels[2] = 10.0;  // 10% jitter
            jitter_levels[3] = 15.0;  // 15% jitter
            
            for (j = 0; j < 4; j = j + 1) begin
                $display("Testing with %.1f%% jitter", jitter_levels[j]);
                
                // Reset and reacquire lock
                rst_n = 0;
                #100;
                rst_n = 1;
                #100;
                
                // Send training with jitter
                for (i = 0; i < 100; i = i + 1) begin
                    send_manchester_bit(i % 2, jitter_levels[j]);
                end
                
                if (locked) begin
                    $display("CDR locked with %.1f%% jitter", jitter_levels[j]);
                end else begin
                    $warning("CDR failed to lock with %.1f%% jitter", jitter_levels[j]);
                end
            end
            
            $display("Jitter tolerance test completed");
        end
    endtask
    
    task bit_error_injection_test;
        integer i;
        integer start_errors;
        begin
            `TEST_SECTION("Bit Error Injection")
            
            // Ensure locked
            if (!locked) begin
                send_training_sequence(100);
                wait(locked);
            end
            
            start_errors = bit_errors;
            
            // Send data with 1% error rate (10000 ppm)
            $display("Sending data with 1%% bit error rate");
            for (i = 0; i < 100; i = i + 1) begin
                send_with_errors(i % 2, 10000);
            end
            
            $display("Bit errors detected: %0d", bit_errors - start_errors);
            
            // CDR should maintain lock despite errors
            `ASSERT(locked === 1'b1, "CDR should maintain lock despite bit errors")
            
            $display("Bit error injection test completed");
        end
    endtask
    
    task lock_maintenance_test;
        integer i;
        integer initial_lock_count;
        begin
            `TEST_SECTION("Lock Maintenance")
            
            // Ensure locked
            if (!locked) begin
                send_training_sequence(100);
                wait(locked);
            end
            
            initial_lock_count = lock_count;
            
            // Send long sequence - lock should be maintained
            $display("Sending 500 bits to test lock maintenance");
            for (i = 0; i < 500; i = i + 1) begin
                send_manchester_bit($random & 1'b1, 0.0);
            end
            
            `ASSERT(locked === 1'b1, "CDR should maintain lock during continuous data")
            `ASSERT(lock_count === initial_lock_count, "Should not lose and reacquire lock")
            
            $display("Lock maintenance test completed");
        end
    endtask
    
    task performance_measurement_test;
        integer start_time, end_time;
        integer num_bits;
        integer start_bits;
        real mbps;
        real ber;
        begin
            `TEST_SECTION("Performance Measurement")
            
            // Ensure locked
            if (!locked) begin
                send_training_sequence(100);
                wait(locked);
            end
            
            num_bits = 200;
            start_time = $time;
            start_bits = bits_received;
            
            // Send random data
            for (integer i = 0; i < num_bits; i = i + 1) begin
                send_manchester_bit($random & 1'b1, 0.0);
            end
            
            end_time = $time;
            
            mbps = (num_bits * 1000.0) / (end_time - start_time);
            ber = (bit_errors * 1.0) / bits_received;
            
            $display("[PERFORMANCE] Recovered %0d bits in %0d ns", 
                     bits_received - start_bits, end_time - start_time);
            $display("[PERFORMANCE] Throughput: %.2f Mbps", mbps);
            $display("[PERFORMANCE] Expected: ~25 Mbps (50 Mbps Manchester / 2)");
            $display("[PERFORMANCE] Bit Error Rate: %.2e", ber);
            $display("[PERFORMANCE] Total lock acquisitions: %0d", lock_count);
            $display("[PERFORMANCE] Total lock losses: %0d", unlock_count);
        end
    endtask

    // ========================================================================
    // Main Test Sequence
    // ========================================================================
    
    initial begin
        // Initialize
        test_failed = 0;
        check_count = 0;
        pass_count = 0;
        fail_count = 0;
        bits_received = 0;
        bit_errors = 0;
        lock_count = 0;
        unlock_count = 0;
        lock_time = 0;
        
        $display("========================================");
        $display("CDR Testbench - Production Grade");
        $display("========================================");
        
        $dumpfile("tb_cdr.vcd");
        $dumpvars(0, tb_cdr);

        // Run test sequence
        reset_test();
        lock_acquisition_test();
        data_recovery_test();
        alternating_pattern_test();
        all_zeros_test();
        all_ones_test();
        jitter_tolerance_test();
        bit_error_injection_test();
        lock_maintenance_test();
        performance_measurement_test();
        
        // Final report
        #1000;
        `TEST_REPORT
        
        $finish;
    end

endmodule
